module top #(
    DATA_WIDTH = 32
) (
    input   logic clk,
    input   logic rst,
    output  logic [DATA_WIDTH-1:0] a0    
);
    
assign a0 = 32'd5;



data_unit1 data_unit(




);












endmodule
