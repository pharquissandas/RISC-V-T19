module pc_pipeline(





);


endmodule
